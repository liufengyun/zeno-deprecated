module Controller (CLK,  busIn, out);
input CLK;
input [31:0] busIn;
output [94:0] out;
wire [3:0] pcNext8;
wire [15:0] instr8;
wire [31:0] stage2Acc8;
wire [146:0] next;
wire out;
reg [51:0] processor8;

assign pcNext8 = ( processor8[51:48] + 4'b0001 );
assign instr8 = ( ( processor8[51:48] == 4'b1111 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1110 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1101 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1100 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1011 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1010 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1001 )? 16'b0000000000000000 : ( ( processor8[51:48] == 4'b1000 )? 16'b0001001100000000 : ( ( processor8[51:48] == 4'b0111 )? 16'b0001000000000010 : ( ( processor8[51:48] == 4'b0110 )? 16'b0000001000000001 : ( ( processor8[51:48] == 4'b0101 )? 16'b0000001001111010 : ( ( processor8[51:48] == 4'b0100 )? 16'b0001000100001000 : ( ( processor8[51:48] == 4'b0011 )? 16'b0000010001111010 : ( ( processor8[51:48] == 4'b0010 )? 16'b0000100100000000 : ( ( processor8[51:48] == 4'b0001 )? 16'b0000100001000001 : ( ( processor8[51:48] == 4'b0000 )? 16'b0000000000000000 : 16'b0000000000000000 ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) );
assign stage2Acc8 = ( ( processor8[15:8] == 8'b00000001 )? ( processor8[47:16] + busIn ) : ( ( processor8[15:8] == 8'b00000011 )? ( processor8[47:16] - busIn ) : ( ( processor8[15:8] == 8'b00000111 )? busIn : ( ( processor8[15:8] == 8'b00001010 )? ( processor8[47:16] & busIn ) : ( ( processor8[15:8] == 8'b00001100 )? ( processor8[47:16] | busIn ) : ( ( processor8[15:8] == 8'b00001110 )? ( ( processor8[47:16] & ~busIn ) | ( ~processor8[47:16] & busIn ) ) : processor8[47:16] ) ) ) ) ) );
assign next = ( ( instr8[15:8] == 8'b00000010 )? {{{pcNext8, ( stage2Acc8 + {24'b000000000000000000000000, instr8[7:0] } ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 + {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000100 )? {{{pcNext8, ( stage2Acc8 - {24'b000000000000000000000000, instr8[7:0] } ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 - {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001000 )? {{{pcNext8, {24'b000000000000000000000000, instr8[7:0] } }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{{24'b000000000000000000000000, instr8[7:0] }, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001001 )? {{{pcNext8, stage2Acc8 }, 16'b0000000000000000 }, {{{{instr8[7:0], 1'b0 }, 1'b1 }, stage2Acc8 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001011 )? {{{pcNext8, ( stage2Acc8 & {24'b000000000000000000000000, instr8[7:0] } ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 & {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001101 )? {{{pcNext8, ( stage2Acc8 | {24'b000000000000000000000000, instr8[7:0] } ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 | {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001111 )? {{{pcNext8, ( ( stage2Acc8 & ~{24'b000000000000000000000000, instr8[7:0] } ) | ( ~stage2Acc8 & {24'b000000000000000000000000, instr8[7:0] } ) ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( ( stage2Acc8 & ~{24'b000000000000000000000000, instr8[7:0] } ) | ( ~stage2Acc8 & {24'b000000000000000000000000, instr8[7:0] } ) ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000101 )? {{{pcNext8, ( stage2Acc8 << instr8[3:0] ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 << instr8[3:0] ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000110 )? {{{pcNext8, ( stage2Acc8 >> instr8[3:0] ) }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( stage2Acc8 >> instr8[3:0] ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010000 )? {{{instr8[3:0], stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, instr8[3:0] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010001 )? ( ( stage2Acc8 == 32'b00000000000000000000000000000000 )? {{{instr8[3:0], stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, instr8[3:0] }, instr8 }, 1'b0 } } } : {{{pcNext8, stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } ) : ( ( instr8[15:8] == 8'b00010010 )? ( ( stage2Acc8 == 32'b00000000000000000000000000000000 )? {{{pcNext8, stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : {{{instr8[3:0], stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, instr8[3:0] }, instr8 }, 1'b0 } } } ) : ( ( instr8[15:8] == 8'b00000001 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000011 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000111 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001010 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001100 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001110 )? {{{pcNext8, stage2Acc8 }, instr8 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010011 )? {{{pcNext8, stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b1 } } } : {{{pcNext8, stage2Acc8 }, 16'b0000000000000000 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{stage2Acc8, pcNext8 }, instr8 }, 1'b0 } } } ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) );
assign out = next[94:0];

initial begin
  processor8 = 52'b0000000000000000000000000000000000000000000000000000;
end

always @ (posedge CLK)
  processor8 <= next[146:95];


endmodule
