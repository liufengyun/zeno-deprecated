module Controller (CLK,  busIn, out);
input CLK;
input [31:0] busIn;
output [96:0] out;
wire [5:0] pcNext8;
wire [15:0] instr8;
wire [135:0] next;
wire [96:0] out;
reg [38:0] processor8;

assign pcNext8 = ( processor8[38:33] + 6'b000001 );
assign instr8 = ( processor8[33]? ( processor8[34]? ( processor8[35]? ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0001000000000010 ) ) ) : ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000010001111010 ) ) ) ) : ( processor8[35]? ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000001001111010 ) ) ) : ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000100001000001 ) ) ) ) ) : ( processor8[34]? ( processor8[35]? ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000001000000001 ) ) ) : ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000100100000000 ) ) ) ) : ( processor8[35]? ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0001000100001000 ) ) ) : ( processor8[36]? ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0001001100000000 ) ) : ( processor8[37]? ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) : ( processor8[38]? 16'b0000000000000000 : 16'b0000000000000000 ) ) ) ) ) );
assign next = ( processor8[0]? ( ( instr8[15:8] == 8'b00000001 )? {{{pcNext8, ( processor8[32:1] + busIn ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] + busIn ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000011 )? {{{pcNext8, ( processor8[32:1] - busIn ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] - busIn ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000111 )? {{{pcNext8, busIn }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{busIn, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001010 )? {{{pcNext8, ( processor8[32:1] & busIn ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] & busIn ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001100 )? {{{pcNext8, ( processor8[32:1] | busIn ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] | busIn ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001110 )? {{{pcNext8, ( ( processor8[32:1] & ~busIn ) | ( ~processor8[32:1] & busIn ) ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( ( processor8[32:1] & ~busIn ) | ( ~processor8[32:1] & busIn ) ), pcNext8 }, instr8 }, 1'b0 } } } : {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b0 } } } ) ) ) ) ) ) : ( ( instr8[15:8] == 8'b00000010 )? {{{pcNext8, ( processor8[32:1] + {24'b000000000000000000000000, instr8[7:0] } ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] + {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000100 )? {{{pcNext8, ( processor8[32:1] - {24'b000000000000000000000000, instr8[7:0] } ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] - {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001000 )? {{{pcNext8, {24'b000000000000000000000000, instr8[7:0] } }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{{24'b000000000000000000000000, instr8[7:0] }, pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001001 )? {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{instr8[7:0], 1'b0 }, 1'b1 }, processor8[32:1] }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001011 )? {{{pcNext8, ( processor8[32:1] & {24'b000000000000000000000000, instr8[7:0] } ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] & {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001101 )? {{{pcNext8, ( processor8[32:1] | {24'b000000000000000000000000, instr8[7:0] } ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] | {24'b000000000000000000000000, instr8[7:0] } ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001111 )? {{{pcNext8, ( ( processor8[32:1] & ~{24'b000000000000000000000000, instr8[7:0] } ) | ( ~processor8[32:1] & {24'b000000000000000000000000, instr8[7:0] } ) ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( ( processor8[32:1] & ~{24'b000000000000000000000000, instr8[7:0] } ) | ( ~processor8[32:1] & {24'b000000000000000000000000, instr8[7:0] } ) ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000101 )? {{{pcNext8, ( processor8[32:1] << instr8[3:0] ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] << instr8[3:0] ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000110 )? {{{pcNext8, ( processor8[32:1] >> instr8[3:0] ) }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{( processor8[32:1] >> instr8[3:0] ), pcNext8 }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010000 )? {{{instr8[5:0], processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], instr8[5:0] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010001 )? ( ( processor8[32:1] == 32'b00000000000000000000000000000000 )? {{{instr8[5:0], processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], instr8[5:0] }, instr8 }, 1'b0 } } } : {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b0 } } } ) : ( ( instr8[15:8] == 8'b00010010 )? ( ( processor8[32:1] == 32'b00000000000000000000000000000000 )? {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b0 } } } : {{{instr8[5:0], processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], instr8[5:0] }, instr8 }, 1'b0 } } } ) : ( ( instr8[15:8] == 8'b00000001 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000011 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00000111 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001010 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001100 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00001110 )? {{{processor8[38:33], processor8[32:1] }, 1'b1 }, {{{{instr8[7:0], 1'b1 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], processor8[38:33] }, instr8 }, 1'b0 } } } : ( ( instr8[15:8] == 8'b00010011 )? {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b1 } } } : {{{pcNext8, processor8[32:1] }, 1'b0 }, {{{{8'b00000000, 1'b0 }, 1'b0 }, 32'b00000000000000000000000000000000 }, {{{processor8[32:1], pcNext8 }, instr8 }, 1'b0 } } } ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) ) );
assign out = next[96:0];

initial begin
  processor8 = 39'b000000000000000000000000000000000000000;
end

always @ (posedge CLK)
  processor8 <= next[135:97];


endmodule
