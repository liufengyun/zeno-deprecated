module Adder ( a, b, out);
input [1:0] a;
input [1:0] b;
output [2:0] out;
wire [2:0] out;


assign out = {{( ( ( ( a[1] & ~b[1] ) | ( ~a[1] & b[1] ) ) & ~( ( x632 & ~1'b0 ) | ( ~( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & 1'b0 ) ) ) | ( ~( ( a[1] & ~b[1] ) | ( ~a[1] & b[1] ) ) & ( ( ( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & ~1'b0 ) | ( ~( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & 1'b0 ) ) ) ), ( ( ( ( a[1] & ~b[1] ) | ( ~a[1] & b[1] ) ) & x591 ) | ( ~( ( a[1] & ~b[1] ) | ( ~a[1] & b[1] ) ) & ( ( ( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & ~1'b0 ) | ( ~( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & 1'b0 ) ) ) ) }, ( ( ( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & ~1'b0 ) | ( ~( ( a[0] & ~b[0] ) | ( ~a[0] & b[0] ) ) & 1'b0 ) ) };


endmodule
